`timescale 1ns/1ns 
module RAM_memory_TB;
	wire [3:0]DataOut;
	reg Enable, ReadWrite,clk;
	reg [3:0]DataIn;
	reg [5:0]Address;
RAM_memory UUT(.Enable(Enable),.ReadWrite(ReadWrite),.clk(clk),.DataIn(DataIn),.Address(Address),.DataOut(DataOut));

initial
	begin
		$dumpfile("RAM_memory.vcd");
		$dumpvars(1,RAM_memory_TB);
			clk=1'b0; #1
			{Enable,ReadWrite,DataIn,Address}=12'b0;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1101010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10000111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10111100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11101010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100011110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101000100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101101111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101110010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110000001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110011110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110101001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111101110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111111110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1001011101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1001100110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1001111001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1010101000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1100000111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1100001101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1100100011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1100110000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10000010101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10001001011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10001101110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10010100010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10100010011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10100100101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10101011011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10110010100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10110110101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10111011101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10111100000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10111110111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11000011011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11010011101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11011111100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100000100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100011001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100110010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100110110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11101010110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11101101001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11111010110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11111100100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11111111001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100000110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100011000110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100011001010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100011100101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100100110111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100101000010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100110100001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100111001111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100111110110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101000001110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101001010110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101001111001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101010111110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101100000110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101100010001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101100110001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101100110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101101010000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101101010100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110000101111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110000111111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110010110001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110100001010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110100110110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110101011100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110101100111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110110001010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110110110001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110110110011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110110111000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110111010011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110111010100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110111110101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110111111111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111000011001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111000100011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111000101001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111000111011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111001001101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111010001011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111010011100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111010101011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111011001000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111011011101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111100001101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111100011010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111100101110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111101110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111110111111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111111001101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111111011110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111111111010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111111111111;#1

		$finish;
	end
	always #1 clk=~clk;
endmodule