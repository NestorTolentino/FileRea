`timescale 1ns/1ns
module mux4_1_TB;
reg [3:0]i1,i2,i3,i4;
reg [1:0]s;
wire [3:0]ot;
mux4_1 UUT(.i2(i2),.i3(i3),.i4(i4),.());
initial
	begin
		$dumpfile("mux4_1.vcd");
		$dumpvars(1,mux4_1_TB);
		{i2,i3,i4}=18'b0;#1
		{i2,i3,i4}=18'b11110011010;#1
		{i2,i3,i4}=18'b100001010100;#1
		{i2,i3,i4}=18'b1110110000010;#1
		{i2,i3,i4}=18'b10101010010111;#1
		{i2,i3,i4}=18'b100101011011100;#1
		{i2,i3,i4}=18'b101110100110010;#1
		{i2,i3,i4}=18'b110000100100101;#1
		{i2,i3,i4}=18'b110001011000010;#1
		{i2,i3,i4}=18'b111100011111110;#1
		{i2,i3,i4}=18'b111110010110000;#1
		{i2,i3,i4}=18'b111110011001101;#1
		{i2,i3,i4}=18'b1000001000111110;#1
		{i2,i3,i4}=18'b1000011000010001;#1
		{i2,i3,i4}=18'b1000100101011101;#1
		{i2,i3,i4}=18'b1000111101010100;#1
		{i2,i3,i4}=18'b1001010001001010;#1
		{i2,i3,i4}=18'b1001100001101001;#1
		{i2,i3,i4}=18'b1001101000110010;#1
		{i2,i3,i4}=18'b1001111010110100;#1
		{i2,i3,i4}=18'b1010010001011100;#1
		{i2,i3,i4}=18'b1100001000110011;#1
		{i2,i3,i4}=18'b1100011001111110;#1
		{i2,i3,i4}=18'b1100110010101111;#1
		{i2,i3,i4}=18'b1100110111100111;#1
		{i2,i3,i4}=18'b1101110001010001;#1
		{i2,i3,i4}=18'b1111100100101110;#1
		{i2,i3,i4}=18'b10001101100011000;#1
		{i2,i3,i4}=18'b10010011111111000;#1
		{i2,i3,i4}=18'b10011000010100011;#1
		{i2,i3,i4}=18'b10100000111110010;#1
		{i2,i3,i4}=18'b10101100001011100;#1
		{i2,i3,i4}=18'b10101100011101100;#1
		{i2,i3,i4}=18'b10101101011101001;#1
		{i2,i3,i4}=18'b10101110011111111;#1
		{i2,i3,i4}=18'b10111001001100011;#1
		{i2,i3,i4}=18'b10111011110010110;#1
		{i2,i3,i4}=18'b11000110100111100;#1
		{i2,i3,i4}=18'b11010001100010111;#1
		{i2,i3,i4}=18'b11011101000110001;#1
		{i2,i3,i4}=18'b11011110100111101;#1
		{i2,i3,i4}=18'b11011110110101011;#1
		{i2,i3,i4}=18'b11110000101000110;#1
		{i2,i3,i4}=18'b11111100001110100;#1
		{i2,i3,i4}=18'b100000011011111011;#1
		{i2,i3,i4}=18'b100000111101110110;#1
		{i2,i3,i4}=18'b100001101001110000;#1
		{i2,i3,i4}=18'b100001111100101001;#1
		{i2,i3,i4}=18'b100010001100011011;#1
		{i2,i3,i4}=18'b100010010101011010;#1
		{i2,i3,i4}=18'b100100100000011010;#1
		{i2,i3,i4}=18'b100100111000101010;#1
		{i2,i3,i4}=18'b100101111100000001;#1
		{i2,i3,i4}=18'b100111011010011011;#1
		{i2,i3,i4}=18'b101000100111101100;#1
		{i2,i3,i4}=18'b101010010000111000;#1
		{i2,i3,i4}=18'b101010100011010100;#1
		{i2,i3,i4}=18'b101010100111100011;#1
		{i2,i3,i4}=18'b101011000100000101;#1
		{i2,i3,i4}=18'b101011101101000011;#1
		{i2,i3,i4}=18'b101100001001000001;#1
		{i2,i3,i4}=18'b101100010000001110;#1
		{i2,i3,i4}=18'b101100100000111110;#1
		{i2,i3,i4}=18'b101101001101101011;#1
		{i2,i3,i4}=18'b101101010000111011;#1
		{i2,i3,i4}=18'b101101011110101011;#1
		{i2,i3,i4}=18'b101101110111101001;#1
		{i2,i3,i4}=18'b101110100111101000;#1
		{i2,i3,i4}=18'b101111000010000111;#1
		{i2,i3,i4}=18'b101111101101100110;#1
		{i2,i3,i4}=18'b110000000001111100;#1
		{i2,i3,i4}=18'b110001111011111011;#1
		{i2,i3,i4}=18'b110010001101100111;#1
		{i2,i3,i4}=18'b110010001111000110;#1
		{i2,i3,i4}=18'b110010010001010100;#1
		{i2,i3,i4}=18'b110100001011101100;#1
		{i2,i3,i4}=18'b110100001110001101;#1
		{i2,i3,i4}=18'b110100010101100111;#1
		{i2,i3,i4}=18'b110100100001110011;#1
		{i2,i3,i4}=18'b110101000000001101;#1
		{i2,i3,i4}=18'b110101100010111010;#1
		{i2,i3,i4}=18'b110111111111011011;#1
		{i2,i3,i4}=18'b111000010001011110;#1
		{i2,i3,i4}=18'b111000011001000001;#1
		{i2,i3,i4}=18'b111000110010110010;#1
		{i2,i3,i4}=18'b111000110111011100;#1
		{i2,i3,i4}=18'b111010100001011000;#1
		{i2,i3,i4}=18'b111010110111111100;#1
		{i2,i3,i4}=18'b111011100111101010;#1
		{i2,i3,i4}=18'b111100010011001001;#1
		{i2,i3,i4}=18'b111101000011001101;#1
		{i2,i3,i4}=18'b111101010010100001;#1
		{i2,i3,i4}=18'b111101011110001111;#1
		{i2,i3,i4}=18'b111101011110011111;#1
		{i2,i3,i4}=18'b111101011110110111;#1
		{i2,i3,i4}=18'b111101100101011010;#1
		{i2,i3,i4}=18'b111110000011000110;#1
		{i2,i3,i4}=18'b111110010001011000;#1
		{i2,i3,i4}=18'b111111010100100001;#1
		{i2,i3,i4}=18'b111111100011100001;#1
		{i2,i3,i4}=18'b111111100100000010;#1
		{i2,i3,i4}=18'b111111111111111111;#1
		$finish;
	end
endmodule
