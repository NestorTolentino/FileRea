`timescale 1ns/1ns 
module RAM_memory_TB;
	wire [3:0]DataOut;
	reg Enable, ReadWrite,clk;
	reg [3:0]DataIn;
	reg [5:0]Address;
RAM_memory UUT(.Enable(Enable),.ReadWrite(ReadWrite),.clk(clk),.DataIn(DataIn),.Address(Address),.DataOut(DataOut));

initial
	begin
		$dumpfile("RAM_memory.vcd");
		$dumpvars(1,RAM_memory_TB);
			clk=1'b0; #1
			{Enable,ReadWrite,DataIn,Address}=12'b0;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1111010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10000010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10110010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11101101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11111101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100000011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100010101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101000101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101001111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101100001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101110111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110001100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111010111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111011010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111011100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1001001001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1001011000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1001111000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1001111101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1010110111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1011111111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1100011101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1100100100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1100101101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1101011111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1101100100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1101100111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1101111001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1110001001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1110011111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1110110001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1110111001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b1111010111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10000010011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10000101010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10001000010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10001101100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10010011100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10011011100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10100111010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10110001010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10110100101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b10111110101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11001001011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11010000001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11010011000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11010110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11011100001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100010010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100101110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11100110010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11101101001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11101111001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11101111100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11110000111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11110010001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11110110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11111100110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11111101000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b11111111010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100000000100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100010000010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100010010000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100011000101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100100101010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100100111010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b100111101001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101000110001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101001100110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101001101111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101010111011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101010111101;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101011010110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101100100100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101101000110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101101110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101110100010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101110101000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b101111111000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110001001000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110001001110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110001011011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110011000111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110011010111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110101000010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110110001011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110110011110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110111010011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b110111110100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111000100001;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111001100100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111001101110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111010100000;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111100010111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111101000010;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111101110110;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111101111111;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111110000011;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111110000100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111110010100;#1
			{Enable,ReadWrite,DataIn,Address}=12'b111111111111;#1

		$finish;
	end
	always #1 clk=~clk;
endmodule