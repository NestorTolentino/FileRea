`timescale 1ns/1ns
module mux4_1_TB;
reg [3:0]i1,i2,i3,i4;
reg [1:0]s;
wire [3:0]ot;
mux4_1 UUT(.i1(i1),.i2(i2),.i3(i3),.i4(i4),.s(s),.ot(ot));
initial
	begin
		$dumpfile("mux4_1.vcd");
		$dumpvars(1,mux4_1_TB);
		{i1,i2,i3,i4,s}=18'b0;#1
		{i1,i2,i3,i4,s}=18'b000000011011001011;#1
		{i1,i2,i3,i4,s}=18'b000000111101100010;#1
		{i1,i2,i3,i4,s}=18'b000001000010010011;#1
		{i1,i2,i3,i4,s}=18'b000001001001101001;#1
		{i1,i2,i3,i4,s}=18'b000001110001101100;#1
		{i1,i2,i3,i4,s}=18'b000001111001011000;#1
		{i1,i2,i3,i4,s}=18'b000010011111010110;#1
		{i1,i2,i3,i4,s}=18'b000010111001011001;#1
		{i1,i2,i3,i4,s}=18'b000011000001011001;#1
		{i1,i2,i3,i4,s}=18'b000100110011000010;#1
		{i1,i2,i3,i4,s}=18'b000101000001001001;#1
		{i1,i2,i3,i4,s}=18'b000110111110110110;#1
		{i1,i2,i3,i4,s}=18'b000111000011000110;#1
		{i1,i2,i3,i4,s}=18'b000111000100100000;#1
		{i1,i2,i3,i4,s}=18'b000111000110100110;#1
		{i1,i2,i3,i4,s}=18'b000111010011111100;#1
		{i1,i2,i3,i4,s}=18'b000111100111111111;#1
		{i1,i2,i3,i4,s}=18'b001001000010100011;#1
		{i1,i2,i3,i4,s}=18'b001001101101100000;#1
		{i1,i2,i3,i4,s}=18'b001010011111010001;#1
		{i1,i2,i3,i4,s}=18'b001011100000011011;#1
		{i1,i2,i3,i4,s}=18'b001011111101011111;#1
		{i1,i2,i3,i4,s}=18'b001100110101011101;#1
		{i1,i2,i3,i4,s}=18'b001101000001001010;#1
		{i1,i2,i3,i4,s}=18'b001101011100110101;#1
		{i1,i2,i3,i4,s}=18'b001101101001010111;#1
		{i1,i2,i3,i4,s}=18'b001110101101001000;#1
		{i1,i2,i3,i4,s}=18'b001111000011011110;#1
		{i1,i2,i3,i4,s}=18'b001111011111010000;#1
		{i1,i2,i3,i4,s}=18'b001111110110110100;#1
		{i1,i2,i3,i4,s}=18'b010001010000010010;#1
		{i1,i2,i3,i4,s}=18'b010001100110000110;#1
		{i1,i2,i3,i4,s}=18'b010001101001001010;#1
		{i1,i2,i3,i4,s}=18'b010010011101001011;#1
		{i1,i2,i3,i4,s}=18'b010011000000000010;#1
		{i1,i2,i3,i4,s}=18'b010101100111011111;#1
		{i1,i2,i3,i4,s}=18'b010110000011101111;#1
		{i1,i2,i3,i4,s}=18'b010110011111011100;#1
		{i1,i2,i3,i4,s}=18'b010111111000000001;#1
		{i1,i2,i3,i4,s}=18'b011000110100001100;#1
		{i1,i2,i3,i4,s}=18'b011001010001111111;#1
		{i1,i2,i3,i4,s}=18'b011010101011111111;#1
		{i1,i2,i3,i4,s}=18'b011011101001100010;#1
		{i1,i2,i3,i4,s}=18'b011101100111100000;#1
		{i1,i2,i3,i4,s}=18'b011110101010100001;#1
		{i1,i2,i3,i4,s}=18'b011111001110001010;#1
		{i1,i2,i3,i4,s}=18'b011111011110110010;#1
		{i1,i2,i3,i4,s}=18'b011111110000100100;#1
		{i1,i2,i3,i4,s}=18'b100000010010010010;#1
		{i1,i2,i3,i4,s}=18'b100001100000110000;#1
		{i1,i2,i3,i4,s}=18'b100001101101110011;#1
		{i1,i2,i3,i4,s}=18'b100010001111001000;#1
		{i1,i2,i3,i4,s}=18'b100010011110000100;#1
		{i1,i2,i3,i4,s}=18'b100100101110001001;#1
		{i1,i2,i3,i4,s}=18'b100100111101110100;#1
		{i1,i2,i3,i4,s}=18'b100101010011010001;#1
		{i1,i2,i3,i4,s}=18'b100101110101101010;#1
		{i1,i2,i3,i4,s}=18'b100111011011001011;#1
		{i1,i2,i3,i4,s}=18'b100111011100111110;#1
		{i1,i2,i3,i4,s}=18'b101000001101000000;#1
		{i1,i2,i3,i4,s}=18'b101000101010011110;#1
		{i1,i2,i3,i4,s}=18'b101001100010101010;#1
		{i1,i2,i3,i4,s}=18'b101001101110001100;#1
		{i1,i2,i3,i4,s}=18'b101001110110100100;#1
		{i1,i2,i3,i4,s}=18'b101001111000111110;#1
		{i1,i2,i3,i4,s}=18'b101010010000101011;#1
		{i1,i2,i3,i4,s}=18'b101010011000110000;#1
		{i1,i2,i3,i4,s}=18'b101011000100101011;#1
		{i1,i2,i3,i4,s}=18'b101011100011011010;#1
		{i1,i2,i3,i4,s}=18'b101011110001101100;#1
		{i1,i2,i3,i4,s}=18'b101011110010010100;#1
		{i1,i2,i3,i4,s}=18'b101011111111001111;#1
		{i1,i2,i3,i4,s}=18'b101100010011100101;#1
		{i1,i2,i3,i4,s}=18'b101100100001001010;#1
		{i1,i2,i3,i4,s}=18'b101100111110111011;#1
		{i1,i2,i3,i4,s}=18'b101101011001011001;#1
		{i1,i2,i3,i4,s}=18'b101101101001001010;#1
		{i1,i2,i3,i4,s}=18'b101111100100011000;#1
		{i1,i2,i3,i4,s}=18'b110001101011001101;#1
		{i1,i2,i3,i4,s}=18'b110100000100011010;#1
		{i1,i2,i3,i4,s}=18'b110100001011111011;#1
		{i1,i2,i3,i4,s}=18'b110100011101010011;#1
		{i1,i2,i3,i4,s}=18'b110110010111111101;#1
		{i1,i2,i3,i4,s}=18'b110111000111000001;#1
		{i1,i2,i3,i4,s}=18'b110111101111100000;#1
		{i1,i2,i3,i4,s}=18'b111000000001001101;#1
		{i1,i2,i3,i4,s}=18'b111000110100011010;#1
		{i1,i2,i3,i4,s}=18'b111010000110010001;#1
		{i1,i2,i3,i4,s}=18'b111011010010001011;#1
		{i1,i2,i3,i4,s}=18'b111011101000011010;#1
		{i1,i2,i3,i4,s}=18'b111011101110001101;#1
		{i1,i2,i3,i4,s}=18'b111011111010000011;#1
		{i1,i2,i3,i4,s}=18'b111100001100000111;#1
		{i1,i2,i3,i4,s}=18'b111100100101011110;#1
		{i1,i2,i3,i4,s}=18'b111100111011010010;#1
		{i1,i2,i3,i4,s}=18'b111101000011010110;#1
		{i1,i2,i3,i4,s}=18'b111110110100010010;#1
		{i1,i2,i3,i4,s}=18'b111111100111001100;#1
		{i1,i2,i3,i4,s}=18'b111111101100001010;#1
		{i1,i2,i3,i4,s}=18'b111111111111111111;#1
		$finish;
	end
endmodule
