`timescale 1ns/1ns
module reg_memory_TB;
reg [4:0] A1,A2,A3;
reg [31:0] WD3;
reg clk,rst,rw;
wire [31:0] RD1,RD2;
reg_memory UUT(.A1(A1),.A2(A2),.A3(A3),.WD3(WD3),.clk(clk),.rst(rst),.rw(rw),.RD1(RD1),.RD2(RD2));
initial
	begin
		$dumpfile("reg_memory.vcd");
		$dumpvars(1,reg_memory_TB);
		clk=1'b0;#1
		rst=1'b1;#1
		rst=1'b0;#1
		{A1,A2,A3,WD3,rw}=50'b0;#1
		{A1,A2,A3,WD3,rw}=50'b10000101100010001100011011;#1
		{A1,A2,A3,WD3,rw}=50'b10100100000001110110000010;#1
		{A1,A2,A3,WD3,rw}=50'b101000001110010001101100111;#1
		{A1,A2,A3,WD3,rw}=50'b1000000100111000011001000001;#1
		{A1,A2,A3,WD3,rw}=50'b1000001101101100010000001110;#1
		{A1,A2,A3,WD3,rw}=50'b1000111011011011110110101011;#1
		{A1,A2,A3,WD3,rw}=50'b1011000000111110000011000110;#1
		{A1,A2,A3,WD3,rw}=50'b1101111011010111001001100011;#1
		{A1,A2,A3,WD3,rw}=50'b10000100111001111100100101110;#1
		{A1,A2,A3,WD3,rw}=50'b10001100100001100110111100111;#1
		{A1,A2,A3,WD3,rw}=50'b10010001000000000100001010100;#1
		{A1,A2,A3,WD3,rw}=50'b10100000011100000111101110110;#1
		{A1,A2,A3,WD3,rw}=50'b10101001111101010010000111000;#1
		{A1,A2,A3,WD3,rw}=50'b11000100110100111011010011011;#1
		{A1,A2,A3,WD3,rw}=50'b11001010010010101110011111111;#1
		{A1,A2,A3,WD3,rw}=50'b11011111011111101011110011111;#1
		{A1,A2,A3,WD3,rw}=50'b11101010011101101010000111011;#1
		{A1,A2,A3,WD3,rw}=50'b11110011111111111010100100001;#1
		{A1,A2,A3,WD3,rw}=50'b11111000101101110100111101000;#1
		{A1,A2,A3,WD3,rw}=50'b100010001000100001101001110000;#1
		{A1,A2,A3,WD3,rw}=50'b100011100011100001111100101001;#1
		{A1,A2,A3,WD3,rw}=50'b100100010000111010100001011000;#1
		{A1,A2,A3,WD3,rw}=50'b100100011000111011100111101010;#1
		{A1,A2,A3,WD3,rw}=50'b100101011100010011000010100011;#1
		{A1,A2,A3,WD3,rw}=50'b100101111001000101110100110010;#1
		{A1,A2,A3,WD3,rw}=50'b101010010010000111110010110000;#1
		{A1,A2,A3,WD3,rw}=50'b101010111010001001010001001010;#1
		{A1,A2,A3,WD3,rw}=50'b101100101010001000011000010001;#1
		{A1,A2,A3,WD3,rw}=50'b101100110110001001101000110010;#1
		{A1,A2,A3,WD3,rw}=50'b101101000111010101101011101001;#1
		{A1,A2,A3,WD3,rw}=50'b101101010100010111011110010110;#1
		{A1,A2,A3,WD3,rw}=50'b101110101100010100000111110010;#1
		{A1,A2,A3,WD3,rw}=50'b110000000001101100100000111110;#1
		{A1,A2,A3,WD3,rw}=50'b110010011110110010001111000110;#1
		{A1,A2,A3,WD3,rw}=50'b110010111111111111100100000010;#1
		{A1,A2,A3,WD3,rw}=50'b110011001110101011000100000101;#1
		{A1,A2,A3,WD3,rw}=50'b110011010100100010010101011010;#1
		{A1,A2,A3,WD3,rw}=50'b111000000001001000001000111110;#1
		{A1,A2,A3,WD3,rw}=50'b111000010000110111111111011011;#1
		{A1,A2,A3,WD3,rw}=50'b111000010101010101100001011100;#1
		{A1,A2,A3,WD3,rw}=50'b111010100101011111100001110100;#1
		{A1,A2,A3,WD3,rw}=50'b111101000110110101100010111010;#1
		{A1,A2,A3,WD3,rw}=50'b111111001011011011101000110001;#1
		{A1,A2,A3,WD3,rw}=50'b1000001100110101100001001000001;#1
		{A1,A2,A3,WD3,rw}=50'b1000001101001111100010011001001;#1
		{A1,A2,A3,WD3,rw}=50'b1000001101101110001111011111011;#1
		{A1,A2,A3,WD3,rw}=50'b1000011000110111101011110110111;#1
		{A1,A2,A3,WD3,rw}=50'b1000011010100111101000011001101;#1
		{A1,A2,A3,WD3,rw}=50'b1000011011011000110000100100101;#1
		{A1,A2,A3,WD3,rw}=50'b1000100000010111010110111111100;#1
		{A1,A2,A3,WD3,rw}=50'b1000101000101101101110111101001;#1
		{A1,A2,A3,WD3,rw}=50'b1000110111010000111110011001101;#1
		{A1,A2,A3,WD3,rw}=50'b1001011010110001000111101010100;#1
		{A1,A2,A3,WD3,rw}=50'b1001101101100010010011111111000;#1
		{A1,A2,A3,WD3,rw}=50'b1001110011010101111101101100110;#1
		{A1,A2,A3,WD3,rw}=50'b1010000011111101101011110101011;#1
		{A1,A2,A3,WD3,rw}=50'b1010001010111110000000001111100;#1
		{A1,A2,A3,WD3,rw}=50'b1010001100110110101000000001101;#1
		{A1,A2,A3,WD3,rw}=50'b1010001111010101101001101101011;#1
		{A1,A2,A3,WD3,rw}=50'b1010100001000101000100111101100;#1
		{A1,A2,A3,WD3,rw}=50'b1010100111001001001111010110100;#1
		{A1,A2,A3,WD3,rw}=50'b1010101011101111111100011100001;#1
		{A1,A2,A3,WD3,rw}=50'b1010111100101000111100011111110;#1
		{A1,A2,A3,WD3,rw}=50'b1010111111001001100110010101111;#1
		{A1,A2,A3,WD3,rw}=50'b1011000000010111101011110001111;#1
		{A1,A2,A3,WD3,rw}=50'b1011011110100000110001011000010;#1
		{A1,A2,A3,WD3,rw}=50'b1011100010010000010101010010111;#1
		{A1,A2,A3,WD3,rw}=50'b1011110100010000100101011011100;#1
		{A1,A2,A3,WD3,rw}=50'b1100001010011111101010010100001;#1
		{A1,A2,A3,WD3,rw}=50'b1100010010101010101100011101100;#1
		{A1,A2,A3,WD3,rw}=50'b1100010100011001000100101011101;#1
		{A1,A2,A3,WD3,rw}=50'b1100010101110111101100101011010;#1
		{A1,A2,A3,WD3,rw}=50'b1100100001111001001100001101001;#1
		{A1,A2,A3,WD3,rw}=50'b1100110001100110100100001110011;#1
		{A1,A2,A3,WD3,rw}=50'b1100110111011110100001110001101;#1
		{A1,A2,A3,WD3,rw}=50'b1100111011000111000010001011110;#1
		{A1,A2,A3,WD3,rw}=50'b1101000010010100100100000011010;#1
		{A1,A2,A3,WD3,rw}=50'b1101010001000110100001011101100;#1
		{A1,A2,A3,WD3,rw}=50'b1101011011010000000011110011010;#1
		{A1,A2,A3,WD3,rw}=50'b1101011100010110100010101100111;#1
		{A1,A2,A3,WD3,rw}=50'b1101100111010101111000010000111;#1
		{A1,A2,A3,WD3,rw}=50'b1101101111010010001101100011000;#1
		{A1,A2,A3,WD3,rw}=50'b1110000101001100100111000101010;#1
		{A1,A2,A3,WD3,rw}=50'b1110001111100110010010001010100;#1
		{A1,A2,A3,WD3,rw}=50'b1110010000111011010001100010111;#1
		{A1,A2,A3,WD3,rw}=50'b1110010010110100000011011111011;#1
		{A1,A2,A3,WD3,rw}=50'b1110011011110111000110111011100;#1
		{A1,A2,A3,WD3,rw}=50'b1110100100110101011101101000011;#1
		{A1,A2,A3,WD3,rw}=50'b1110100101100001101110001010001;#1
		{A1,A2,A3,WD3,rw}=50'b1110101010001011110000101000110;#1
		{A1,A2,A3,WD3,rw}=50'b1110101101000101010100011010100;#1
		{A1,A2,A3,WD3,rw}=50'b1110110010001001010010001011100;#1
		{A1,A2,A3,WD3,rw}=50'b1110111001001001100011001111110;#1
		{A1,A2,A3,WD3,rw}=50'b1110111010001100101111100000001;#1
		{A1,A2,A3,WD3,rw}=50'b1111001100000111000110010110010;#1
		{A1,A2,A3,WD3,rw}=50'b1111001111000101010100111100011;#1
		{A1,A2,A3,WD3,rw}=50'b1111010011011011000110100111100;#1
		{A1,A2,A3,WD3,rw}=50'b1111100001111011011110100111101;#1
		{A1,A2,A3,WD3,rw}=50'b1111100100000111110010001011000;#1
		{A1,A2,A3,WD3,rw}=50'b1111111110111001100001000110011;#1
		{A1,A2,A3,WD3,rw}=50'b11111111111111111111111111111111111111111111111111;#1
		$finish;
	end
	always #1 clk=~clk;
endmodule
