`timescale 1ns/1ns 
module mux4_1_TB;
	wire [3:0]ot;
	reg [3:0]i1,i2,i3,i4;
	reg [1:0]s;
mux4_1 UUT(.i1(i1),.i2(i2),.i3(i3),.i4(i4),.s(s),.ot(ot));

initial
	begin
		$dumpfile("mux4_1.vcd");
		$dumpvars(1,mux4_1_TB);
			{i1,i2,i3,i4,s}=18'b000000000000000000;#1
			{i1,i2,i3,i4,s}=18'b111110000111100101;#1
			{i1,i2,i3,i4,s}=18'b011101101000110011;#1
			{i1,i2,i3,i4,s}=18'b110101000100110100;#1
			{i1,i2,i3,i4,s}=18'b000101000010111001;#1
			{i1,i2,i3,i4,s}=18'b010110100101100011;#1
			{i1,i2,i3,i4,s}=18'b100101000010000111;#1
			{i1,i2,i3,i4,s}=18'b000101010111100111;#1
			{i1,i2,i3,i4,s}=18'b100101000000100100;#1
			{i1,i2,i3,i4,s}=18'b001101111001110111;#1
			{i1,i2,i3,i4,s}=18'b110100010011011111;#1
			{i1,i2,i3,i4,s}=18'b101001001111010100;#1
			{i1,i2,i3,i4,s}=18'b101010100101111101;#1
			{i1,i2,i3,i4,s}=18'b110000001100001010;#1
			{i1,i2,i3,i4,s}=18'b011101000010001100;#1
			{i1,i2,i3,i4,s}=18'b011011101010110111;#1
			{i1,i2,i3,i4,s}=18'b111010111111000110;#1
			{i1,i2,i3,i4,s}=18'b101011111011110001;#1
			{i1,i2,i3,i4,s}=18'b111110000011100011;#1
			{i1,i2,i3,i4,s}=18'b101100001100001010;#1
			{i1,i2,i3,i4,s}=18'b000100111000101000;#1
			{i1,i2,i3,i4,s}=18'b011000000101101011;#1
			{i1,i2,i3,i4,s}=18'b101010111100001010;#1
			{i1,i2,i3,i4,s}=18'b100001001001011000;#1
			{i1,i2,i3,i4,s}=18'b111110111000001100;#1
			{i1,i2,i3,i4,s}=18'b101110011001001110;#1
			{i1,i2,i3,i4,s}=18'b111101010111111011;#1
			{i1,i2,i3,i4,s}=18'b101001111011011001;#1
			{i1,i2,i3,i4,s}=18'b001101001100011011;#1
			{i1,i2,i3,i4,s}=18'b111110011001000010;#1
			{i1,i2,i3,i4,s}=18'b100100000110110110;#1
			{i1,i2,i3,i4,s}=18'b000000100100000100;#1
			{i1,i2,i3,i4,s}=18'b011111001000111010;#1
			{i1,i2,i3,i4,s}=18'b111101110010010010;#1
			{i1,i2,i3,i4,s}=18'b000111100101011110;#1
			{i1,i2,i3,i4,s}=18'b001100100010101010;#1
			{i1,i2,i3,i4,s}=18'b100110000000011110;#1
			{i1,i2,i3,i4,s}=18'b001111100010000001;#1
			{i1,i2,i3,i4,s}=18'b110000011010101101;#1
			{i1,i2,i3,i4,s}=18'b110000111000001110;#1
			{i1,i2,i3,i4,s}=18'b101011011111000111;#1
			{i1,i2,i3,i4,s}=18'b110011010000101111;#1
			{i1,i2,i3,i4,s}=18'b000001001101011010;#1
			{i1,i2,i3,i4,s}=18'b100011010100000100;#1
			{i1,i2,i3,i4,s}=18'b001101010000110010;#1
			{i1,i2,i3,i4,s}=18'b000001001001000111;#1
			{i1,i2,i3,i4,s}=18'b101100110010111011;#1
			{i1,i2,i3,i4,s}=18'b010010101100011000;#1
			{i1,i2,i3,i4,s}=18'b100000011100101011;#1
			{i1,i2,i3,i4,s}=18'b000101011010101000;#1
			{i1,i2,i3,i4,s}=18'b111110111111011101;#1
			{i1,i2,i3,i4,s}=18'b001101101110111100;#1
			{i1,i2,i3,i4,s}=18'b010011011110010111;#1
			{i1,i2,i3,i4,s}=18'b101100100100100111;#1
			{i1,i2,i3,i4,s}=18'b010001000010110000;#1
			{i1,i2,i3,i4,s}=18'b010111100010110000;#1
			{i1,i2,i3,i4,s}=18'b111000100111111010;#1
			{i1,i2,i3,i4,s}=18'b010110111000000011;#1
			{i1,i2,i3,i4,s}=18'b100101110011011000;#1
			{i1,i2,i3,i4,s}=18'b011000010000101110;#1
			{i1,i2,i3,i4,s}=18'b110100100101110110;#1
			{i1,i2,i3,i4,s}=18'b001011000100000001;#1
			{i1,i2,i3,i4,s}=18'b000111110100100011;#1
			{i1,i2,i3,i4,s}=18'b000101100001100111;#1
			{i1,i2,i3,i4,s}=18'b010010000010010100;#1
			{i1,i2,i3,i4,s}=18'b001011010011110010;#1
			{i1,i2,i3,i4,s}=18'b110100000111111100;#1
			{i1,i2,i3,i4,s}=18'b110010100100110100;#1
			{i1,i2,i3,i4,s}=18'b010101001110010001;#1
			{i1,i2,i3,i4,s}=18'b011101000101000100;#1
			{i1,i2,i3,i4,s}=18'b101000011001100101;#1
			{i1,i2,i3,i4,s}=18'b110110101101000101;#1
			{i1,i2,i3,i4,s}=18'b111001000000000110;#1
			{i1,i2,i3,i4,s}=18'b111001000000000101;#1
			{i1,i2,i3,i4,s}=18'b000000011100110010;#1
			{i1,i2,i3,i4,s}=18'b011100001011101110;#1
			{i1,i2,i3,i4,s}=18'b000101110000010101;#1
			{i1,i2,i3,i4,s}=18'b110110001110100110;#1
			{i1,i2,i3,i4,s}=18'b011000110000110110;#1
			{i1,i2,i3,i4,s}=18'b101011000001001111;#1
			{i1,i2,i3,i4,s}=18'b010001010000110110;#1
			{i1,i2,i3,i4,s}=18'b110001001011010001;#1
			{i1,i2,i3,i4,s}=18'b110111111110111001;#1
			{i1,i2,i3,i4,s}=18'b001101110101011111;#1
			{i1,i2,i3,i4,s}=18'b000000111111111011;#1
			{i1,i2,i3,i4,s}=18'b011001000110001100;#1
			{i1,i2,i3,i4,s}=18'b001011000101001101;#1
			{i1,i2,i3,i4,s}=18'b101001000101110100;#1
			{i1,i2,i3,i4,s}=18'b011110011110111001;#1
			{i1,i2,i3,i4,s}=18'b000010010001010001;#1
			{i1,i2,i3,i4,s}=18'b110101010100010100;#1
			{i1,i2,i3,i4,s}=18'b011111110101001110;#1
			{i1,i2,i3,i4,s}=18'b111100001010101110;#1
			{i1,i2,i3,i4,s}=18'b100011001101110000;#1
			{i1,i2,i3,i4,s}=18'b010111101101101101;#1
			{i1,i2,i3,i4,s}=18'b101100011101010100;#1
			{i1,i2,i3,i4,s}=18'b000100000101001111;#1
			{i1,i2,i3,i4,s}=18'b100100100100000011;#1
			{i1,i2,i3,i4,s}=18'b111011111000111011;#1
			{i1,i2,i3,i4,s}=18'b011000011110000110;#1
			{i1,i2,i3,i4,s}=18'b001101101001011001;#1
			{i1,i2,i3,i4,s}=18'b111111111111111111;#1

		$finish;
	end

endmodule